-- example from: https://jnjsite.com/vhdl-sumador-completo-de-1-bit/
-- Sumador completo de 1 bit

-- Librerías

library IEEE;
use IEEE.std_logic_1164.all;


-- Declaración de la entidad del circuito

entity oneBitFullAdder is
    port (
        sum, carryOut : out std_logic;
        a, b, carryIn : in std_logic
    );
end entity;

-- Arquitectura del circuito

architecture arch of oneBitFullAdder is
begin

    sum <= ((not carryIn) and (not a) and b)
        or ((not carryIn) and a and (not b))
        or (carryIn and (not a) and (not b))
        or (carryIn and a and b);

    carryOut <= (carryIn and b) or (a and b) or (carryIn and a);

end architecture;
