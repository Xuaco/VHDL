-- example from: https://jnjsite.com/vhdl-sumador-completo-de-1-bit/
-- Sumador completo de 1 bit

-- Librerías



-- Declaración de la entidad del circuito



-- Arquitectura del circuito
